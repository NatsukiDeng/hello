module moduleName (
);
    
    wire one;

endmodule