module moduleName (
);
    
    //push this
    //mod

endmodule