module moduleName (
);
    
    //push this

endmodule